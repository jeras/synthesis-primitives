///////////////////////////////////////////////////////////////////////////////
// Extended Golay encoder,
// testbench
//
// Copyright 2025 Iztok Jeras <iztok.jeras@gmail.com>
//
// Licensed under CERN-OHL-P v2 or later
///////////////////////////////////////////////////////////////////////////////

import golay_pkg::*;

module golay_tb();

endmodule: golay_tb;