module crash ();

    localparam logic [4-1:0] max_lst [5] = '{0, 1, 2**4-1};

endmodule: crash
