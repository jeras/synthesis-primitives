///////////////////////////////////////////////////////////////////////////////
// Extended Golay code package
//
// Copyright 2025 Iztok Jeras <iztok.jeras@gmail.com>
//
// Licensed under CERN-OHL-P v2 or later
///////////////////////////////////////////////////////////////////////////////

package golay_pkg;

    logic [0:24-1] golay_matrix [0:12-1] = '{
        24'b100000000000_100111110001,
        24'b010000000000_010011111010,
        24'b001000000000_001001111101,
        24'b000100000000_100100111110,
        24'b000010000000_110010011101,
        24'b000001000000_111001001110,
        24'b000000100000_111100100101,
        24'b000000010000_111110010010,
        24'b000000001000_011111001001,
        24'b000000000100_001111100110,
        24'b000000000010_010101010111,
        24'b000000000001_101010101011
    };

endpackage: golay_pkg
